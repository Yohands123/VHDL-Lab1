LIBRARY ieee; 
USE ieee.std_logic_1164.all; 
LIBRARY work; 
ENTITY VHDL_Polarity_Controller IS
	PORT(
		POLARITY_CONTROL, IN_1, IN_2, IN_3, IN_4 : IN STD_LOGIC; 
		OUT_1, OUT_2, OUT_3, OUT_4 : OUT STD_LOGIC
		); 

END ENTITY VHDL_Polarity_Controller; 


ARCHITECTURE polarity_control OF VHDL_Polarity_Controller IS
BEGIN

OUT_1 <= POLARITY_CONTROL XNOR IN_1;
OUT_2 <= POLARITY_CONTROL XNOR IN_2;
OUT_3 <= POLARITY_CONTROL XNOR IN_3;
OUT_4 <= POLARITY_CONTROL XNOR IN_4;

END polarity_control; 